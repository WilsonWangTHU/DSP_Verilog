library verilog;
use verilog.vl_types.all;
entity LED_FLOW is
end LED_FLOW;
