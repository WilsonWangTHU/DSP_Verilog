library verilog;
use verilog.vl_types.all;
entity test_encode_decode_outof_module is
end test_encode_decode_outof_module;
