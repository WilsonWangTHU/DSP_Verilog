library verilog;
use verilog.vl_types.all;
entity test_encode_decode is
end test_encode_decode;
