library verilog;
use verilog.vl_types.all;
entity test_ask is
end test_ask;
